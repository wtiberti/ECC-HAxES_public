-- Component: tb_FullAdder
-- Desc: Testbed for the FullAdder component
-- Author: Walter Tiberti <walter.tiberti@graduate.univaq.it>

library ieee;
use ieee.std_logic_1164.all;

entity tb_FullAdder is
end tb_FullAdder;

architecture rtl of tb_FullAdder is

begin

end rtl;
